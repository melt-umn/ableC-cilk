grammar edu:umn:cs:melt:exts:ableC:cilk:src:concretesyntax;

exports edu:umn:cs:melt:exts:ableC:cilk:src:concretesyntax:functionDef;
exports edu:umn:cs:melt:exts:ableC:cilk:src:concretesyntax:returnStmt;
exports edu:umn:cs:melt:exts:ableC:cilk:src:concretesyntax:syncStmt;
exports edu:umn:cs:melt:exts:ableC:cilk:src:concretesyntax:spawnExpr;
exports edu:umn:cs:melt:exts:ableC:cilk:src:concretesyntax:exitStmt;


