grammar edu:umn:cs:melt:exts:ableC:cilk:src ;

exports edu:umn:cs:melt:exts:ableC:cilk:src:abstractsyntax ;
exports edu:umn:cs:melt:exts:ableC:cilk:src:concretesyntax ;

