grammar edu:umn:cs:melt:exts:ableC:cilk:concretesyntax;

import edu:umn:cs:melt:ableC:concretesyntax;

marking terminal Cilk_t 'cilk' lexer classes {Ckeyword};
