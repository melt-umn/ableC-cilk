grammar edu:umn:cs:melt:exts:ableC:cilk:src:concretesyntax;

exports edu:umn:cs:melt:exts:ableC:cilk:src:concretesyntax:cilk;
exports edu:umn:cs:melt:exts:ableC:cilk:src:concretesyntax:syncStmt;
exports edu:umn:cs:melt:exts:ableC:cilk:src:concretesyntax:spawnStmt;
exports edu:umn:cs:melt:exts:ableC:cilk:src:concretesyntax:exitStmt;


