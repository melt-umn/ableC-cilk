grammar edu:umn:cs:melt:exts:ableC:cilk;

exports edu:umn:cs:melt:exts:ableC:cilk:abstractsyntax;
exports edu:umn:cs:melt:exts:ableC:cilk:concretesyntax;

