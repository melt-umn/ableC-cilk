grammar edu:umn:cs:melt:exts:ableC:cilk:abstractsyntax; 

imports silver:langutil;
imports silver:langutil:pp with implode as ppImplode, concat as ppConcat;
