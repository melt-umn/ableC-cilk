grammar edu:umn:cs:melt:exts:ableC:cilk:concretesyntax;

exports edu:umn:cs:melt:exts:ableC:cilk:concretesyntax:functionDef;
exports edu:umn:cs:melt:exts:ableC:cilk:concretesyntax:returnStmt;
exports edu:umn:cs:melt:exts:ableC:cilk:concretesyntax:syncStmt;
exports edu:umn:cs:melt:exts:ableC:cilk:concretesyntax:spawnStmt;
exports edu:umn:cs:melt:exts:ableC:cilk:concretesyntax:exitStmt;


